localparam CHAR_CR = 8'h0D;
localparam CHAR_LF = 8'h0A;

localparam CHAR_SP = 8'h20;

localparam CHAR_0 = 8'h30;
localparam CHAR_1 = 8'h31;
localparam CHAR_2 = 8'h32;
localparam CHAR_3 = 8'h33;
localparam CHAR_4 = 8'h34;
localparam CHAR_5 = 8'h35;
localparam CHAR_6 = 8'h36;
localparam CHAR_7 = 8'h37;
localparam CHAR_8 = 8'h38;
localparam CHAR_9 = 8'h39;

localparam CHAR_QM = 8'h3F;

localparam CHAR_A = 8'h41;
localparam CHAR_B = 8'h42;
localparam CHAR_C = 8'h43;
localparam CHAR_D = 8'h44;
localparam CHAR_E = 8'h45;
localparam CHAR_F = 8'h46;
localparam CHAR_G = 8'h47;
localparam CHAR_H = 8'h48;
localparam CHAR_I = 8'h49;
localparam CHAR_J = 8'h4A;
localparam CHAR_K = 8'h4B;
localparam CHAR_L = 8'h4C;
localparam CHAR_M = 8'h4D;
localparam CHAR_N = 8'h4E;
localparam CHAR_O = 8'h4F;
localparam CHAR_P = 8'h50;
localparam CHAR_Q = 8'h51;
localparam CHAR_R = 8'h52;
localparam CHAR_S = 8'h53;
localparam CHAR_T = 8'h54;
localparam CHAR_U = 8'h55;
localparam CHAR_V = 8'h56;
localparam CHAR_W = 8'h57;
localparam CHAR_X = 8'h58;
localparam CHAR_Y = 8'h59;
localparam CHAR_Z = 8'h5A;

localparam CHAR_a = 8'h61;
localparam CHAR_b = 8'h62;
localparam CHAR_c = 8'h63;
localparam CHAR_d = 8'h64;
localparam CHAR_e = 8'h65;
localparam CHAR_f = 8'h66;
localparam CHAR_g = 8'h67;
localparam CHAR_h = 8'h68;
localparam CHAR_i = 8'h69;
localparam CHAR_j = 8'h6A;
localparam CHAR_k = 8'h6B;
localparam CHAR_l = 8'h6C;
localparam CHAR_m = 8'h6D;
localparam CHAR_n = 8'h6E;
localparam CHAR_o = 8'h6F;
localparam CHAR_p = 8'h70;
localparam CHAR_q = 8'h71;
localparam CHAR_r = 8'h72;
localparam CHAR_s = 8'h73;
localparam CHAR_t = 8'h74;
localparam CHAR_u = 8'h75;
localparam CHAR_v = 8'h76;
localparam CHAR_w = 8'h77;
localparam CHAR_x = 8'h78;
localparam CHAR_y = 8'h79;
localparam CHAR_z = 8'h7A;
