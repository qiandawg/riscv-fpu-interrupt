/************************************************
  The Verilog HDL code example is from the book
  Computer Principles and Design in Verilog HDL
  by Yamin Li, published by A JOHN WILEY & SONS
************************************************/
module wallace_26x24 (a,b,x,y,z);                      // 26*24 wallace tree
    input  [25:00] b;                                  // 26 bits
    input  [23:00] a;                                  // 24 bits
    output [49:08] x;                                  // sum high
    output [49:08] y;                                  // carry high
    output [07:00] z;                                  // sum low
    reg    [25:00] p [23:00];                          // p[i][j]
    parameter zero = 1'b0;                             // constant 0
    integer i, j;
    always @ * begin
        for (i = 0; i < 24; i = i + 1)
            for (j = 0; j < 26; j = j + 1)
                p[i][j] = a[i] & b[j];                 // p[i][j]=a[i]&b[j]
    end
    // level 1 ------------------------------------------------------------
    wire  [7:0] s1 [46:1];
    wire  [7:0] c1 [47:2];
    //     49:
    //     48:   p[23][25]
    //     47:   p[22][25], p[23][24]
    csa a1_46_0 (p[21][25], p[22][24], p[23][23], s1[46][0], c1[47][0]);
    csa a1_45_0 (p[20][25], p[21][24], p[22][23], s1[45][0], c1[46][0]);
    //     45:   p[23][22]
    csa a1_44_1 (p[19][25], p[20][24], p[21][23], s1[44][1], c1[45][1]);
    csa a1_44_0 (p[22][22], p[23][21],      zero, s1[44][0], c1[45][0]);
    csa a1_43_1 (p[18][25], p[19][24], p[20][23], s1[43][1], c1[44][1]);
    csa a1_43_0 (p[21][22], p[22][21], p[23][20], s1[43][0], c1[44][0]);
    csa a1_42_1 (p[17][25], p[18][24], p[19][23], s1[42][1], c1[43][1]);
    csa a1_42_0 (p[20][22], p[21][21], p[22][20], s1[42][0], c1[43][0]);
    //     42:   p[23][19]
    csa a1_41_2 (p[16][25], p[17][24], p[18][23], s1[41][2], c1[42][2]);
    csa a1_41_1 (p[19][22], p[20][21], p[21][20], s1[41][1], c1[42][1]);
    csa a1_41_0 (p[22][19], p[23][18],      zero, s1[41][0], c1[42][0]);
    csa a1_40_2 (p[15][25], p[16][24], p[17][23], s1[40][2], c1[41][2]);
    csa a1_40_1 (p[18][22], p[19][21], p[20][20], s1[40][1], c1[41][1]);
    csa a1_40_0 (p[21][19], p[22][18], p[23][17], s1[40][0], c1[41][0]);
    csa a1_39_2 (p[14][25], p[15][24], p[16][23], s1[39][2], c1[40][2]);
    csa a1_39_1 (p[17][22], p[18][21], p[19][20], s1[39][1], c1[40][1]);
    csa a1_39_0 (p[20][19], p[21][18], p[22][17], s1[39][0], c1[40][0]);
    //     39:   p[23][16]
    csa a1_38_3 (p[13][25], p[14][24], p[15][23], s1[38][3], c1[39][3]);
    csa a1_38_2 (p[16][22], p[17][21], p[18][20], s1[38][2], c1[39][2]);
    csa a1_38_1 (p[19][19], p[20][18], p[21][17], s1[38][1], c1[39][1]);
    csa a1_38_0 (p[22][16], p[23][15],      zero, s1[38][0], c1[39][0]);
    csa a1_37_3 (p[12][25], p[13][24], p[14][23], s1[37][3], c1[38][3]);
    csa a1_37_2 (p[15][22], p[16][21], p[17][20], s1[37][2], c1[38][2]);
    csa a1_37_1 (p[18][19], p[19][18], p[20][17], s1[37][1], c1[38][1]);
    csa a1_37_0 (p[21][16], p[22][15], p[23][14], s1[37][0], c1[38][0]);
    csa a1_36_3 (p[11][25], p[12][24], p[13][23], s1[36][3], c1[37][3]);
    csa a1_36_2 (p[14][22], p[15][21], p[16][20], s1[36][2], c1[37][2]);
    csa a1_36_1 (p[17][19], p[18][18], p[19][17], s1[36][1], c1[37][1]);
    csa a1_36_0 (p[20][16], p[21][15], p[22][14], s1[36][0], c1[37][0]);
    //     36:   p[23][13]
    csa a1_35_4 (p[10][25], p[11][24], p[12][23], s1[35][4], c1[36][4]);
    csa a1_35_3 (p[13][22], p[14][21], p[15][20], s1[35][3], c1[36][3]);
    csa a1_35_2 (p[16][19], p[17][18], p[18][17], s1[35][2], c1[36][2]);
    csa a1_35_1 (p[19][16], p[20][15], p[21][14], s1[35][1], c1[36][1]);
    csa a1_35_0 (p[22][13], p[23][12],      zero, s1[35][0], c1[36][0]);
    csa a1_34_4 (p[09][25], p[10][24], p[11][23], s1[34][4], c1[35][4]);
    csa a1_34_3 (p[12][22], p[13][21], p[14][20], s1[34][3], c1[35][3]);
    csa a1_34_2 (p[15][19], p[16][18], p[17][17], s1[34][2], c1[35][2]);
    csa a1_34_1 (p[18][16], p[19][15], p[20][14], s1[34][1], c1[35][1]);
    csa a1_34_0 (p[21][13], p[22][12], p[23][11], s1[34][0], c1[35][0]);
    csa a1_33_4 (p[08][25], p[09][24], p[10][23], s1[33][4], c1[34][4]);
    csa a1_33_3 (p[11][22], p[12][21], p[13][20], s1[33][3], c1[34][3]);
    csa a1_33_2 (p[14][19], p[15][18], p[16][17], s1[33][2], c1[34][2]);
    csa a1_33_1 (p[17][16], p[18][15], p[19][14], s1[33][1], c1[34][1]);
    csa a1_33_0 (p[20][13], p[21][12], p[22][11], s1[33][0], c1[34][0]);
    //     33:   p[23][10]
    csa a1_32_5 (p[07][25], p[08][24], p[09][23], s1[32][5], c1[33][5]);
    csa a1_32_4 (p[10][22], p[11][21], p[12][20], s1[32][4], c1[33][4]);
    csa a1_32_3 (p[13][19], p[14][18], p[15][17], s1[32][3], c1[33][3]);
    csa a1_32_2 (p[16][16], p[17][15], p[18][14], s1[32][2], c1[33][2]);
    csa a1_32_1 (p[19][13], p[20][12], p[21][11], s1[32][1], c1[33][1]);
    csa a1_32_0 (p[22][10], p[23][09],      zero, s1[32][0], c1[33][0]);
    csa a1_31_5 (p[06][25], p[07][24], p[08][23], s1[31][5], c1[32][5]);
    csa a1_31_4 (p[09][22], p[10][21], p[11][20], s1[31][4], c1[32][4]);
    csa a1_31_3 (p[12][19], p[13][18], p[14][17], s1[31][3], c1[32][3]);
    csa a1_31_2 (p[15][16], p[16][15], p[17][14], s1[31][2], c1[32][2]);
    csa a1_31_1 (p[18][13], p[19][12], p[20][11], s1[31][1], c1[32][1]);
    csa a1_31_0 (p[21][10], p[22][09], p[23][08], s1[31][0], c1[32][0]);
    csa a1_30_5 (p[05][25], p[06][24], p[07][23], s1[30][5], c1[31][5]);
    csa a1_30_4 (p[08][22], p[09][21], p[10][20], s1[30][4], c1[31][4]);
    csa a1_30_3 (p[11][19], p[12][18], p[13][17], s1[30][3], c1[31][3]);
    csa a1_30_2 (p[14][16], p[15][15], p[16][14], s1[30][2], c1[31][2]);
    csa a1_30_1 (p[17][13], p[18][12], p[19][11], s1[30][1], c1[31][1]);
    csa a1_30_0 (p[20][10], p[21][09], p[22][08], s1[30][0], c1[31][0]);
    //     30:   p[23][07]
    csa a1_29_6 (p[04][25], p[05][24], p[06][23], s1[29][6], c1[30][6]);
    csa a1_29_5 (p[07][22], p[08][21], p[09][20], s1[29][5], c1[30][5]);
    csa a1_29_4 (p[10][19], p[11][18], p[12][17], s1[29][4], c1[30][4]);
    csa a1_29_3 (p[13][16], p[14][15], p[15][14], s1[29][3], c1[30][3]);
    csa a1_29_2 (p[16][13], p[17][12], p[18][11], s1[29][2], c1[30][2]);
    csa a1_29_1 (p[19][10], p[20][09], p[21][08], s1[29][1], c1[30][1]);
    csa a1_29_0 (p[22][07], p[23][06],      zero, s1[29][0], c1[30][0]);
    csa a1_28_6 (p[03][25], p[04][24], p[05][23], s1[28][6], c1[29][6]);
    csa a1_28_5 (p[06][22], p[07][21], p[08][20], s1[28][5], c1[29][5]);
    csa a1_28_4 (p[09][19], p[10][18], p[11][17], s1[28][4], c1[29][4]);
    csa a1_28_3 (p[12][16], p[13][15], p[14][14], s1[28][3], c1[29][3]);
    csa a1_28_2 (p[15][13], p[16][12], p[17][11], s1[28][2], c1[29][2]);
    csa a1_28_1 (p[18][10], p[19][09], p[20][08], s1[28][1], c1[29][1]);
    csa a1_28_0 (p[21][07], p[22][06], p[23][05], s1[28][0], c1[29][0]);
    csa a1_27_6 (p[02][25], p[03][24], p[04][23], s1[27][6], c1[28][6]);
    csa a1_27_5 (p[05][22], p[06][21], p[07][20], s1[27][5], c1[28][5]);
    csa a1_27_4 (p[08][19], p[09][18], p[10][17], s1[27][4], c1[28][4]);
    csa a1_27_3 (p[11][16], p[12][15], p[13][14], s1[27][3], c1[28][3]);
    csa a1_27_2 (p[14][13], p[15][12], p[16][11], s1[27][2], c1[28][2]);
    csa a1_27_1 (p[17][10], p[18][09], p[19][08], s1[27][1], c1[28][1]);
    csa a1_27_0 (p[20][07], p[21][06], p[22][05], s1[27][0], c1[28][0]);
    //     27:   p[23][04]
    csa a1_26_7 (p[01][25], p[02][24], p[03][23], s1[26][7], c1[27][7]);
    csa a1_26_6 (p[04][22], p[05][21], p[06][20], s1[26][6], c1[27][6]);
    csa a1_26_5 (p[07][19], p[08][18], p[09][17], s1[26][5], c1[27][5]);
    csa a1_26_4 (p[10][16], p[11][15], p[12][14], s1[26][4], c1[27][4]);
    csa a1_26_3 (p[13][13], p[14][12], p[15][11], s1[26][3], c1[27][3]);
    csa a1_26_2 (p[16][10], p[17][09], p[18][08], s1[26][2], c1[27][2]);
    csa a1_26_1 (p[19][07], p[20][06], p[21][05], s1[26][1], c1[27][1]);
    csa a1_26_0 (p[22][04], p[23][03],      zero, s1[26][0], c1[27][0]);
    csa a1_25_7 (p[00][25], p[01][24], p[02][23], s1[25][7], c1[26][7]);
    csa a1_25_6 (p[03][22], p[04][21], p[05][20], s1[25][6], c1[26][6]);
    csa a1_25_5 (p[06][19], p[07][18], p[08][17], s1[25][5], c1[26][5]);
    csa a1_25_4 (p[09][16], p[10][15], p[11][14], s1[25][4], c1[26][4]);
    csa a1_25_3 (p[12][13], p[13][12], p[14][11], s1[25][3], c1[26][3]);
    csa a1_25_2 (p[15][10], p[16][09], p[17][08], s1[25][2], c1[26][2]);
    csa a1_25_1 (p[18][07], p[19][06], p[20][05], s1[25][1], c1[26][1]);
    csa a1_25_0 (p[21][04], p[22][03], p[23][02], s1[25][0], c1[26][0]);
    csa a1_24_7 (p[00][24], p[01][23], p[02][22], s1[24][7], c1[25][7]);
    csa a1_24_6 (p[03][21], p[04][20], p[05][19], s1[24][6], c1[25][6]);
    csa a1_24_5 (p[06][18], p[07][17], p[08][16], s1[24][5], c1[25][5]);
    csa a1_24_4 (p[09][15], p[10][14], p[11][13], s1[24][4], c1[25][4]);
    csa a1_24_3 (p[12][12], p[13][11], p[14][10], s1[24][3], c1[25][3]);
    csa a1_24_2 (p[15][09], p[16][08], p[17][07], s1[24][2], c1[25][2]);
    csa a1_24_1 (p[18][06], p[19][05], p[20][04], s1[24][1], c1[25][1]);
    csa a1_24_0 (p[21][03], p[22][02], p[23][01], s1[24][0], c1[25][0]);
    csa a1_23_7 (p[00][23], p[01][22], p[02][21], s1[23][7], c1[24][7]);
    csa a1_23_6 (p[03][20], p[04][19], p[05][18], s1[23][6], c1[24][6]);
    csa a1_23_5 (p[06][17], p[07][16], p[08][15], s1[23][5], c1[24][5]);
    csa a1_23_4 (p[09][14], p[10][13], p[11][12], s1[23][4], c1[24][4]);
    csa a1_23_3 (p[12][11], p[13][10], p[14][09], s1[23][3], c1[24][3]);
    csa a1_23_2 (p[15][08], p[16][07], p[17][06], s1[23][2], c1[24][2]);
    csa a1_23_1 (p[18][05], p[19][04], p[20][03], s1[23][1], c1[24][1]);
    csa a1_23_0 (p[21][02], p[22][01], p[23][00], s1[23][0], c1[24][0]);
    csa a1_22_7 (p[00][22], p[01][21], p[02][20], s1[22][7], c1[23][7]);
    csa a1_22_6 (p[03][19], p[04][18], p[05][17], s1[22][6], c1[23][6]);
    csa a1_22_5 (p[06][16], p[07][15], p[08][14], s1[22][5], c1[23][5]);
    csa a1_22_4 (p[09][13], p[10][12], p[11][11], s1[22][4], c1[23][4]);
    csa a1_22_3 (p[12][10], p[13][09], p[14][08], s1[22][3], c1[23][3]);
    csa a1_22_2 (p[15][07], p[16][06], p[17][05], s1[22][2], c1[23][2]);
    csa a1_22_1 (p[18][04], p[19][03], p[20][02], s1[22][1], c1[23][1]);
    csa a1_22_0 (p[21][01], p[22][00],      zero, s1[22][0], c1[23][0]);
    csa a1_21_6 (p[00][21], p[01][20], p[02][19], s1[21][6], c1[22][6]);
    csa a1_21_5 (p[03][18], p[04][17], p[05][16], s1[21][5], c1[22][5]);
    csa a1_21_4 (p[06][15], p[07][14], p[08][13], s1[21][4], c1[22][4]);
    csa a1_21_3 (p[09][12], p[10][11], p[11][10], s1[21][3], c1[22][3]);
    csa a1_21_2 (p[12][09], p[13][08], p[14][07], s1[21][2], c1[22][2]);
    csa a1_21_1 (p[15][06], p[16][05], p[17][04], s1[21][1], c1[22][1]);
    csa a1_21_0 (p[18][03], p[19][02], p[20][01], s1[21][0], c1[22][0]);
    //     21:   p[21][00]
    csa a1_20_6 (p[00][20], p[01][19], p[02][18], s1[20][6], c1[21][6]);
    csa a1_20_5 (p[03][17], p[04][16], p[05][15], s1[20][5], c1[21][5]);
    csa a1_20_4 (p[06][14], p[07][13], p[08][12], s1[20][4], c1[21][4]);
    csa a1_20_3 (p[09][11], p[10][10], p[11][09], s1[20][3], c1[21][3]);
    csa a1_20_2 (p[12][08], p[13][07], p[14][06], s1[20][2], c1[21][2]);
    csa a1_20_1 (p[15][05], p[16][04], p[17][03], s1[20][1], c1[21][1]);
    csa a1_20_0 (p[18][02], p[19][01], p[20][00], s1[20][0], c1[21][0]);
    csa a1_19_6 (p[00][19], p[01][18], p[02][17], s1[19][6], c1[20][6]);
    csa a1_19_5 (p[03][16], p[04][15], p[05][14], s1[19][5], c1[20][5]);
    csa a1_19_4 (p[06][13], p[07][12], p[08][11], s1[19][4], c1[20][4]);
    csa a1_19_3 (p[09][10], p[10][09], p[11][08], s1[19][3], c1[20][3]);
    csa a1_19_2 (p[12][07], p[13][06], p[14][05], s1[19][2], c1[20][2]);
    csa a1_19_1 (p[15][04], p[16][03], p[17][02], s1[19][1], c1[20][1]);
    csa a1_19_0 (p[18][01], p[19][00],      zero, s1[19][0], c1[20][0]);
    csa a1_18_5 (p[00][18], p[01][17], p[02][16], s1[18][5], c1[19][5]);
    csa a1_18_4 (p[03][15], p[04][14], p[05][13], s1[18][4], c1[19][4]);
    csa a1_18_3 (p[06][12], p[07][11], p[08][10], s1[18][3], c1[19][3]);
    csa a1_18_2 (p[09][09], p[10][08], p[11][07], s1[18][2], c1[19][2]);
    csa a1_18_1 (p[12][06], p[13][05], p[14][04], s1[18][1], c1[19][1]);
    csa a1_18_0 (p[15][03], p[16][02], p[17][01], s1[18][0], c1[19][0]);
    //     18:   p[18][00]
    csa a1_17_5 (p[00][17], p[01][16], p[02][15], s1[17][5], c1[18][5]);
    csa a1_17_4 (p[03][14], p[04][13], p[05][12], s1[17][4], c1[18][4]);
    csa a1_17_3 (p[06][11], p[07][10], p[08][09], s1[17][3], c1[18][3]);
    csa a1_17_2 (p[09][08], p[10][07], p[11][06], s1[17][2], c1[18][2]);
    csa a1_17_1 (p[12][05], p[13][04], p[14][03], s1[17][1], c1[18][1]);
    csa a1_17_0 (p[15][02], p[16][01], p[17][00], s1[17][0], c1[18][0]);
    csa a1_16_5 (p[00][16], p[01][15], p[02][14], s1[16][5], c1[17][5]);
    csa a1_16_4 (p[03][13], p[04][12], p[05][11], s1[16][4], c1[17][4]);
    csa a1_16_3 (p[06][10], p[07][09], p[08][08], s1[16][3], c1[17][3]);
    csa a1_16_2 (p[09][07], p[10][06], p[11][05], s1[16][2], c1[17][2]);
    csa a1_16_1 (p[12][04], p[13][03], p[14][02], s1[16][1], c1[17][1]);
    csa a1_16_0 (p[15][01], p[16][00],      zero, s1[16][0], c1[17][0]);
    csa a1_15_4 (p[00][15], p[01][14], p[02][13], s1[15][4], c1[16][4]);
    csa a1_15_3 (p[03][12], p[04][11], p[05][10], s1[15][3], c1[16][3]);
    csa a1_15_2 (p[06][09], p[07][08], p[08][07], s1[15][2], c1[16][2]);
    csa a1_15_1 (p[09][06], p[10][05], p[11][04], s1[15][1], c1[16][1]);
    csa a1_15_0 (p[12][03], p[13][02], p[14][01], s1[15][0], c1[16][0]);
    //     15:   p[15][00]
    csa a1_14_4 (p[00][14], p[01][13], p[02][12], s1[14][4], c1[15][4]);
    csa a1_14_3 (p[03][11], p[04][10], p[05][09], s1[14][3], c1[15][3]);
    csa a1_14_2 (p[06][08], p[07][07], p[08][06], s1[14][2], c1[15][2]);
    csa a1_14_1 (p[09][05], p[10][04], p[11][03], s1[14][1], c1[15][1]);
    csa a1_14_0 (p[12][02], p[13][01], p[14][00], s1[14][0], c1[15][0]);
    csa a1_13_4 (p[00][13], p[01][12], p[02][11], s1[13][4], c1[14][4]);
    csa a1_13_3 (p[03][10], p[04][09], p[05][08], s1[13][3], c1[14][3]);
    csa a1_13_2 (p[06][07], p[07][06], p[08][05], s1[13][2], c1[14][2]);
    csa a1_13_1 (p[09][04], p[10][03], p[11][02], s1[13][1], c1[14][1]);
    csa a1_13_0 (p[12][01], p[13][00],      zero, s1[13][0], c1[14][0]);
    csa a1_12_3 (p[00][12], p[01][11], p[02][10], s1[12][3], c1[13][3]);
    csa a1_12_2 (p[03][09], p[04][08], p[05][07], s1[12][2], c1[13][2]);
    csa a1_12_1 (p[06][06], p[07][05], p[08][04], s1[12][1], c1[13][1]);
    csa a1_12_0 (p[09][03], p[10][02], p[11][01], s1[12][0], c1[13][0]);
    //     12:   p[12][00]
    csa a1_11_3 (p[00][11], p[01][10], p[02][09], s1[11][3], c1[12][3]);
    csa a1_11_2 (p[03][08], p[04][07], p[05][06], s1[11][2], c1[12][2]);
    csa a1_11_1 (p[06][05], p[07][04], p[08][03], s1[11][1], c1[12][1]);
    csa a1_11_0 (p[09][02], p[10][01], p[11][00], s1[11][0], c1[12][0]);
    csa a1_10_3 (p[00][10], p[01][09], p[02][08], s1[10][3], c1[11][3]);
    csa a1_10_2 (p[03][07], p[04][06], p[05][05], s1[10][2], c1[11][2]);
    csa a1_10_1 (p[06][04], p[07][03], p[08][02], s1[10][1], c1[11][1]);
    csa a1_10_0 (p[09][01], p[10][00],      zero, s1[10][0], c1[11][0]);
    csa a1_09_2 (p[00][09], p[01][08], p[02][07], s1[09][2], c1[10][2]);
    csa a1_09_1 (p[03][06], p[04][05], p[05][04], s1[09][1], c1[10][1]);
    csa a1_09_0 (p[06][03], p[07][02], p[08][01], s1[09][0], c1[10][0]);
    //     09:   p[09][00]
    csa a1_08_2 (p[00][08], p[01][07], p[02][06], s1[08][2], c1[09][2]);
    csa a1_08_1 (p[03][05], p[04][04], p[05][03], s1[08][1], c1[09][1]);
    csa a1_08_0 (p[06][02], p[07][01], p[08][00], s1[08][0], c1[09][0]);
    csa a1_07_2 (p[00][07], p[01][06], p[02][05], s1[07][2], c1[08][2]);
    csa a1_07_1 (p[03][04], p[04][03], p[05][02], s1[07][1], c1[08][1]);
    csa a1_07_0 (p[06][01], p[07][00],      zero, s1[07][0], c1[08][0]);
    csa a1_06_1 (p[00][06], p[01][05], p[02][04], s1[06][1], c1[07][1]);
    csa a1_06_0 (p[03][03], p[04][02], p[05][01], s1[06][0], c1[07][0]);
    //     06:   p[06][00]
    csa a1_05_1 (p[00][05], p[01][04], p[02][03], s1[05][1], c1[06][1]);
    csa a1_05_0 (p[03][02], p[04][01], p[05][00], s1[05][0], c1[06][0]);
    csa a1_04_1 (p[00][04], p[01][03], p[02][02], s1[04][1], c1[05][1]);
    csa a1_04_0 (p[03][01], p[04][00],      zero, s1[04][0], c1[05][0]);
    csa a1_03_0 (p[00][03], p[01][02], p[02][01], s1[03][0], c1[04][0]);
    //     03:   p[03][00]
    csa a1_02_0 (p[00][02], p[01][01], p[02][00], s1[02][0], c1[03][0]);
    csa a1_01_0 (p[00][01], p[01][00],      zero, s1[01][0], c1[02][0]);
    //     00:   p[00][00]
    // level 2 ------------------------------------------------------------
    wire  [4:0] s2 [47:2];
    wire  [4:0] c2 [48:3];
    //     49:
    //     48:   p[23][25]
    csa a2_47_0 (p[22][25], p[23][24], c1[47][0], s2[47][0], c2[48][0]);
    csa a2_46_0 (s1[46][0], c1[46][0],      zero, s2[46][0], c2[47][0]);
    csa a2_45_0 (s1[45][0], p[23][22], c1[45][1], s2[45][0], c2[46][0]);
    //     45:   c1[45][0]
    csa a2_44_0 (s1[44][1], s1[44][0], c1[44][1], s2[44][0], c2[45][0]);
    //     44:   c1[44][0]
    csa a2_43_0 (s1[43][1], s1[43][0], c1[43][1], s2[43][0], c2[44][0]);
    //     43:   c1[43][0]
    csa a2_42_1 (s1[42][1], s1[42][0], p[23][19], s2[42][1], c2[43][1]);
    csa a2_42_0 (c1[42][2], c1[42][1], c1[42][0], s2[42][0], c2[43][0]);
    csa a2_41_1 (s1[41][2], s1[41][1], s1[41][0], s2[41][1], c2[42][1]);
    csa a2_41_0 (c1[41][2], c1[41][1], c1[41][0], s2[41][0], c2[42][0]);
    csa a2_40_1 (s1[40][2], s1[40][1], s1[40][0], s2[40][1], c2[41][1]);
    csa a2_40_0 (c1[40][2], c1[40][1], c1[40][0], s2[40][0], c2[41][0]);
    csa a2_39_2 (s1[39][2], s1[39][1], s1[39][0], s2[39][2], c2[40][2]);
    csa a2_39_1 (p[23][16], c1[39][3], c1[39][2], s2[39][1], c2[40][1]);
    csa a2_39_0 (c1[39][1], c1[39][0],      zero, s2[39][0], c2[40][0]);
    csa a2_38_2 (s1[38][3], s1[38][2], s1[38][1], s2[38][2], c2[39][2]);
    csa a2_38_1 (s1[38][0], c1[38][3], c1[38][2], s2[38][1], c2[39][1]);
    csa a2_38_0 (c1[38][1], c1[38][0],      zero, s2[38][0], c2[39][0]);
    csa a2_37_2 (s1[37][3], s1[37][2], s1[37][1], s2[37][2], c2[38][2]);
    csa a2_37_1 (s1[37][0], c1[37][3], c1[37][2], s2[37][1], c2[38][1]);
    csa a2_37_0 (c1[37][1], c1[37][0],      zero, s2[37][0], c2[38][0]);
    csa a2_36_2 (s1[36][3], s1[36][2], s1[36][1], s2[36][2], c2[37][2]);
    csa a2_36_1 (s1[36][0], p[23][13], c1[36][4], s2[36][1], c2[37][1]);
    csa a2_36_0 (c1[36][3], c1[36][2], c1[36][1], s2[36][0], c2[37][0]);
    //     36:   c1[36][0]
    csa a2_35_2 (s1[35][4], s1[35][3], s1[35][2], s2[35][2], c2[36][2]);
    csa a2_35_1 (s1[35][1], s1[35][0], c1[35][4], s2[35][1], c2[36][1]);
    csa a2_35_0 (c1[35][3], c1[35][2], c1[35][1], s2[35][0], c2[36][0]);
    //     35:   c1[35][0]
    csa a2_34_2 (s1[34][4], s1[34][3], s1[34][2], s2[34][2], c2[35][2]);
    csa a2_34_1 (s1[34][1], s1[34][0], c1[34][4], s2[34][1], c2[35][1]);
    csa a2_34_0 (c1[34][3], c1[34][2], c1[34][1], s2[34][0], c2[35][0]);
    //     34:   c1[34][0]
    csa a2_33_3 (s1[33][4], s1[33][3], s1[33][2], s2[33][3], c2[34][3]);
    csa a2_33_2 (s1[33][1], s1[33][0], p[23][10], s2[33][2], c2[34][2]);
    csa a2_33_1 (c1[33][5], c1[33][4], c1[33][3], s2[33][1], c2[34][1]);
    csa a2_33_0 (c1[33][2], c1[33][1], c1[33][0], s2[33][0], c2[34][0]);
    csa a2_32_3 (s1[32][5], s1[32][4], s1[32][3], s2[32][3], c2[33][3]);
    csa a2_32_2 (s1[32][2], s1[32][1], s1[32][0], s2[32][2], c2[33][2]);
    csa a2_32_1 (c1[32][5], c1[32][4], c1[32][3], s2[32][1], c2[33][1]);
    csa a2_32_0 (c1[32][2], c1[32][1], c1[32][0], s2[32][0], c2[33][0]);
    csa a2_31_3 (s1[31][5], s1[31][4], s1[31][3], s2[31][3], c2[32][3]);
    csa a2_31_2 (s1[31][2], s1[31][1], s1[31][0], s2[31][2], c2[32][2]);
    csa a2_31_1 (c1[31][5], c1[31][4], c1[31][3], s2[31][1], c2[32][1]);
    csa a2_31_0 (c1[31][2], c1[31][1], c1[31][0], s2[31][0], c2[32][0]);
    csa a2_30_4 (s1[30][5], s1[30][4], s1[30][3], s2[30][4], c2[31][4]);
    csa a2_30_3 (s1[30][2], s1[30][1], s1[30][0], s2[30][3], c2[31][3]);
    csa a2_30_2 (p[23][07], c1[30][6], c1[30][5], s2[30][2], c2[31][2]);
    csa a2_30_1 (c1[30][4], c1[30][3], c1[30][2], s2[30][1], c2[31][1]);
    csa a2_30_0 (c1[30][1], c1[30][0],      zero, s2[30][0], c2[31][0]);
    csa a2_29_4 (s1[29][6], s1[29][5], s1[29][4], s2[29][4], c2[30][4]);
    csa a2_29_3 (s1[29][3], s1[29][2], s1[29][1], s2[29][3], c2[30][3]);
    csa a2_29_2 (s1[29][0], c1[29][6], c1[29][5], s2[29][2], c2[30][2]);
    csa a2_29_1 (c1[29][4], c1[29][3], c1[29][2], s2[29][1], c2[30][1]);
    csa a2_29_0 (c1[29][1], c1[29][0],      zero, s2[29][0], c2[30][0]);
    csa a2_28_4 (s1[28][6], s1[28][5], s1[28][4], s2[28][4], c2[29][4]);
    csa a2_28_3 (s1[28][3], s1[28][2], s1[28][1], s2[28][3], c2[29][3]);
    csa a2_28_2 (s1[28][0], c1[28][6], c1[28][5], s2[28][2], c2[29][2]);
    csa a2_28_1 (c1[28][4], c1[28][3], c1[28][2], s2[28][1], c2[29][1]);
    csa a2_28_0 (c1[28][1], c1[28][0],      zero, s2[28][0], c2[29][0]);
    csa a2_27_4 (s1[27][6], s1[27][5], s1[27][4], s2[27][4], c2[28][4]);
    csa a2_27_3 (s1[27][3], s1[27][2], s1[27][1], s2[27][3], c2[28][3]);
    csa a2_27_2 (s1[27][0], p[23][04], c1[27][7], s2[27][2], c2[28][2]);
    csa a2_27_1 (c1[27][6], c1[27][5], c1[27][4], s2[27][1], c2[28][1]);
    csa a2_27_0 (c1[27][3], c1[27][2], c1[27][1], s2[27][0], c2[28][0]);
    //     27:   c1[27][0]
    csa a2_26_4 (s1[26][7], s1[26][6], s1[26][5], s2[26][4], c2[27][4]);
    csa a2_26_3 (s1[26][4], s1[26][3], s1[26][2], s2[26][3], c2[27][3]);
    csa a2_26_2 (s1[26][1], s1[26][0], c1[26][7], s2[26][2], c2[27][2]);
    csa a2_26_1 (c1[26][6], c1[26][5], c1[26][4], s2[26][1], c2[27][1]);
    csa a2_26_0 (c1[26][3], c1[26][2], c1[26][1], s2[26][0], c2[27][0]);
    //     26:   c1[26][0]
    csa a2_25_4 (s1[25][7], s1[25][6], s1[25][5], s2[25][4], c2[26][4]);
    csa a2_25_3 (s1[25][4], s1[25][3], s1[25][2], s2[25][3], c2[26][3]);
    csa a2_25_2 (s1[25][1], s1[25][0], c1[25][7], s2[25][2], c2[26][2]);
    csa a2_25_1 (c1[25][6], c1[25][5], c1[25][4], s2[25][1], c2[26][1]);
    csa a2_25_0 (c1[25][3], c1[25][2], c1[25][1], s2[25][0], c2[26][0]);
    //     25:   c1[25][0]
    csa a2_24_4 (s1[24][7], s1[24][6], s1[24][5], s2[24][4], c2[25][4]);
    csa a2_24_3 (s1[24][4], s1[24][3], s1[24][2], s2[24][3], c2[25][3]);
    csa a2_24_2 (s1[24][1], s1[24][0], c1[24][7], s2[24][2], c2[25][2]);
    csa a2_24_1 (c1[24][6], c1[24][5], c1[24][4], s2[24][1], c2[25][1]);
    csa a2_24_0 (c1[24][3], c1[24][2], c1[24][1], s2[24][0], c2[25][0]);
    //     24:   c1[24][0]
    csa a2_23_4 (s1[23][7], s1[23][6], s1[23][5], s2[23][4], c2[24][4]);
    csa a2_23_3 (s1[23][4], s1[23][3], s1[23][2], s2[23][3], c2[24][3]);
    csa a2_23_2 (s1[23][1], s1[23][0], c1[23][7], s2[23][2], c2[24][2]);
    csa a2_23_1 (c1[23][6], c1[23][5], c1[23][4], s2[23][1], c2[24][1]);
    csa a2_23_0 (c1[23][3], c1[23][2], c1[23][1], s2[23][0], c2[24][0]);
    //     23:   c1[23][0]
    csa a2_22_4 (s1[22][7], s1[22][6], s1[22][5], s2[22][4], c2[23][4]);
    csa a2_22_3 (s1[22][4], s1[22][3], s1[22][2], s2[22][3], c2[23][3]);
    csa a2_22_2 (s1[22][1], s1[22][0], c1[22][6], s2[22][2], c2[23][2]);
    csa a2_22_1 (c1[22][5], c1[22][4], c1[22][3], s2[22][1], c2[23][1]);
    csa a2_22_0 (c1[22][2], c1[22][1], c1[22][0], s2[22][0], c2[23][0]);
    csa a2_21_4 (s1[21][6], s1[21][5], s1[21][4], s2[21][4], c2[22][4]);
    csa a2_21_3 (s1[21][3], s1[21][2], s1[21][1], s2[21][3], c2[22][3]);
    csa a2_21_2 (s1[21][0], p[21][00], c1[21][6], s2[21][2], c2[22][2]);
    csa a2_21_1 (c1[21][5], c1[21][4], c1[21][3], s2[21][1], c2[22][1]);
    csa a2_21_0 (c1[21][2], c1[21][1], c1[21][0], s2[21][0], c2[22][0]);
    csa a2_20_4 (s1[20][6], s1[20][5], s1[20][4], s2[20][4], c2[21][4]);
    csa a2_20_3 (s1[20][3], s1[20][2], s1[20][1], s2[20][3], c2[21][3]);
    csa a2_20_2 (s1[20][0], c1[20][6], c1[20][5], s2[20][2], c2[21][2]);
    csa a2_20_1 (c1[20][4], c1[20][3], c1[20][2], s2[20][1], c2[21][1]);
    csa a2_20_0 (c1[20][1], c1[20][0],      zero, s2[20][0], c2[21][0]);
    csa a2_19_3 (s1[19][6], s1[19][5], s1[19][4], s2[19][3], c2[20][3]);
    csa a2_19_2 (s1[19][3], s1[19][2], s1[19][1], s2[19][2], c2[20][2]);
    csa a2_19_1 (s1[19][0], c1[19][5], c1[19][4], s2[19][1], c2[20][1]);
    csa a2_19_0 (c1[19][3], c1[19][2], c1[19][1], s2[19][0], c2[20][0]);
    //     19:   c1[19][0]
    csa a2_18_3 (s1[18][5], s1[18][4], s1[18][3], s2[18][3], c2[19][3]);
    csa a2_18_2 (s1[18][2], s1[18][1], s1[18][0], s2[18][2], c2[19][2]);
    csa a2_18_1 (p[18][00], c1[18][5], c1[18][4], s2[18][1], c2[19][1]);
    csa a2_18_0 (c1[18][3], c1[18][2], c1[18][1], s2[18][0], c2[19][0]);
    //     18:   c1[18][0]
    csa a2_17_3 (s1[17][5], s1[17][4], s1[17][3], s2[17][3], c2[18][3]);
    csa a2_17_2 (s1[17][2], s1[17][1], s1[17][0], s2[17][2], c2[18][2]);
    csa a2_17_1 (c1[17][5], c1[17][4], c1[17][3], s2[17][1], c2[18][1]);
    csa a2_17_0 (c1[17][2], c1[17][1], c1[17][0], s2[17][0], c2[18][0]);
    csa a2_16_3 (s1[16][5], s1[16][4], s1[16][3], s2[16][3], c2[17][3]);
    csa a2_16_2 (s1[16][2], s1[16][1], s1[16][0], s2[16][2], c2[17][2]);
    csa a2_16_1 (c1[16][4], c1[16][3], c1[16][2], s2[16][1], c2[17][1]);
    csa a2_16_0 (c1[16][1], c1[16][0],      zero, s2[16][0], c2[17][0]);
    csa a2_15_3 (s1[15][4], s1[15][3], s1[15][2], s2[15][3], c2[16][3]);
    csa a2_15_2 (s1[15][1], s1[15][0], p[15][00], s2[15][2], c2[16][2]);
    csa a2_15_1 (c1[15][4], c1[15][3], c1[15][2], s2[15][1], c2[16][1]);
    csa a2_15_0 (c1[15][1], c1[15][0],      zero, s2[15][0], c2[16][0]);
    csa a2_14_2 (s1[14][4], s1[14][3], s1[14][2], s2[14][2], c2[15][2]);
    csa a2_14_1 (s1[14][1], s1[14][0], c1[14][4], s2[14][1], c2[15][1]);
    csa a2_14_0 (c1[14][3], c1[14][2], c1[14][1], s2[14][0], c2[15][0]);
    //     14:   c1[14][0]
    csa a2_13_2 (s1[13][4], s1[13][3], s1[13][2], s2[13][2], c2[14][2]);
    csa a2_13_1 (s1[13][1], s1[13][0], c1[13][3], s2[13][1], c2[14][1]);
    csa a2_13_0 (c1[13][2], c1[13][1], c1[13][0], s2[13][0], c2[14][0]);
    csa a2_12_2 (s1[12][3], s1[12][2], s1[12][1], s2[12][2], c2[13][2]);
    csa a2_12_1 (s1[12][0], p[12][00], c1[12][3], s2[12][1], c2[13][1]);
    csa a2_12_0 (c1[12][2], c1[12][1], c1[12][0], s2[12][0], c2[13][0]);
    csa a2_11_2 (s1[11][3], s1[11][2], s1[11][1], s2[11][2], c2[12][2]);
    csa a2_11_1 (s1[11][0], c1[11][3], c1[11][2], s2[11][1], c2[12][1]);
    csa a2_11_0 (c1[11][1], c1[11][0],      zero, s2[11][0], c2[12][0]);
    csa a2_10_1 (s1[10][3], s1[10][2], s1[10][1], s2[10][1], c2[11][1]);
    csa a2_10_0 (s1[10][0], c1[10][2], c1[10][1], s2[10][0], c2[11][0]);
    //     10:   c1[10][0]
    csa a2_09_1 (s1[09][2], s1[09][1], s1[09][0], s2[09][1], c2[10][1]);
    csa a2_09_0 (p[09][00], c1[09][2], c1[09][1], s2[09][0], c2[10][0]);
    //     09:   c1[09][0]
    csa a2_08_1 (s1[08][2], s1[08][1], s1[08][0], s2[08][1], c2[09][1]);
    csa a2_08_0 (c1[08][2], c1[08][1], c1[08][0], s2[08][0], c2[09][0]);
    csa a2_07_1 (s1[07][2], s1[07][1], s1[07][0], s2[07][1], c2[08][1]);
    csa a2_07_0 (c1[07][1], c1[07][0],      zero, s2[07][0], c2[08][0]);
    csa a2_06_1 (s1[06][1], s1[06][0], p[06][00], s2[06][1], c2[07][1]);
    csa a2_06_0 (c1[06][1], c1[06][0],      zero, s2[06][0], c2[07][0]);
    csa a2_05_0 (s1[05][1], s1[05][0], c1[05][1], s2[05][0], c2[06][0]);
    //     05:   c1[05][0]
    csa a2_04_0 (s1[04][1], s1[04][0], c1[04][0], s2[04][0], c2[05][0]);
    csa a2_03_0 (s1[03][0], p[03][00], c1[03][0], s2[03][0], c2[04][0]);
    csa a2_02_0 (s1[02][0], c1[02][0],      zero, s2[02][0], c2[03][0]);
    //     01:   s1[01][0]
    //     00:   p[00][00]
    // level 3 ------------------------------------------------------------
    wire  [3:0] s3 [48:3];
    wire  [3:0] c3 [49:4];
    //     49:
    csa a3_48_0 (p[23][25], c2[48][0],      zero, s3[48][0], c3[49][0]);
    csa a3_47_0 (s2[47][0], c2[47][0],      zero, s3[47][0], c3[48][0]);
    csa a3_46_0 (s2[46][0], c2[46][0],      zero, s3[46][0], c3[47][0]);
    csa a3_45_0 (s2[45][0], c1[45][0], c2[45][0], s3[45][0], c3[46][0]);
    csa a3_44_0 (s2[44][0], c1[44][0], c2[44][0], s3[44][0], c3[45][0]);
    csa a3_43_0 (s2[43][0], c1[43][0], c2[43][1], s3[43][0], c3[44][0]);
    //     43:   c2[43][0]
    csa a3_42_0 (s2[42][1], s2[42][0], c2[42][1], s3[42][0], c3[43][0]);
    //     42:   c2[42][0]
    csa a3_41_0 (s2[41][1], s2[41][0], c2[41][1], s3[41][0], c3[42][0]);
    //     41:   c2[41][0]
    csa a3_40_1 (s2[40][1], s2[40][0], c2[40][2], s3[40][1], c3[41][1]);
    csa a3_40_0 (c2[40][1], c2[40][0],      zero, s3[40][0], c3[41][0]);
    csa a3_39_1 (s2[39][2], s2[39][1], s2[39][0], s3[39][1], c3[40][1]);
    csa a3_39_0 (c2[39][2], c2[39][1], c2[39][0], s3[39][0], c3[40][0]);
    csa a3_38_1 (s2[38][2], s2[38][1], s2[38][0], s3[38][1], c3[39][1]);
    csa a3_38_0 (c2[38][2], c2[38][1], c2[38][0], s3[38][0], c3[39][0]);
    csa a3_37_1 (s2[37][2], s2[37][1], s2[37][0], s3[37][1], c3[38][1]);
    csa a3_37_0 (c2[37][2], c2[37][1], c2[37][0], s3[37][0], c3[38][0]);
    csa a3_36_1 (s2[36][2], s2[36][1], s2[36][0], s3[36][1], c3[37][1]);
    csa a3_36_0 (c1[36][0], c2[36][2], c2[36][1], s3[36][0], c3[37][0]);
    //     36:   c2[36][0]
    csa a3_35_1 (s2[35][2], s2[35][1], s2[35][0], s3[35][1], c3[36][1]);
    csa a3_35_0 (c1[35][0], c2[35][2], c2[35][1], s3[35][0], c3[36][0]);
    //     35:   c2[35][0]
    csa a3_34_2 (s2[34][2], s2[34][1], s2[34][0], s3[34][2], c3[35][2]);
    csa a3_34_1 (c1[34][0], c2[34][3], c2[34][2], s3[34][1], c3[35][1]);
    csa a3_34_0 (c2[34][1], c2[34][0],      zero, s3[34][0], c3[35][0]);
    csa a3_33_2 (s2[33][3], s2[33][2], s2[33][1], s3[33][2], c3[34][2]);
    csa a3_33_1 (s2[33][0], c2[33][3], c2[33][2], s3[33][1], c3[34][1]);
    csa a3_33_0 (c2[33][1], c2[33][0],      zero, s3[33][0], c3[34][0]);
    csa a3_32_2 (s2[32][3], s2[32][2], s2[32][1], s3[32][2], c3[33][2]);
    csa a3_32_1 (s2[32][0], c2[32][3], c2[32][2], s3[32][1], c3[33][1]);
    csa a3_32_0 (c2[32][1], c2[32][0],      zero, s3[32][0], c3[33][0]);
    csa a3_31_2 (s2[31][3], s2[31][2], s2[31][1], s3[31][2], c3[32][2]);
    csa a3_31_1 (s2[31][0], c2[31][4], c2[31][3], s3[31][1], c3[32][1]);
    csa a3_31_0 (c2[31][2], c2[31][1], c2[31][0], s3[31][0], c3[32][0]);
    csa a3_30_2 (s2[30][4], s2[30][3], s2[30][2], s3[30][2], c3[31][2]);
    csa a3_30_1 (s2[30][1], s2[30][0], c2[30][4], s3[30][1], c3[31][1]);
    csa a3_30_0 (c2[30][3], c2[30][2], c2[30][1], s3[30][0], c3[31][0]);
    //     30:   c2[30][0]
    csa a3_29_2 (s2[29][4], s2[29][3], s2[29][2], s3[29][2], c3[30][2]);
    csa a3_29_1 (s2[29][1], s2[29][0], c2[29][4], s3[29][1], c3[30][1]);
    csa a3_29_0 (c2[29][3], c2[29][2], c2[29][1], s3[29][0], c3[30][0]);
    //     29:   c2[29][0]
    csa a3_28_2 (s2[28][4], s2[28][3], s2[28][2], s3[28][2], c3[29][2]);
    csa a3_28_1 (s2[28][1], s2[28][0], c2[28][4], s3[28][1], c3[29][1]);
    csa a3_28_0 (c2[28][3], c2[28][2], c2[28][1], s3[28][0], c3[29][0]);
    //     28:   c2[28][0]
    csa a3_27_3 (s2[27][4], s2[27][3], s2[27][2], s3[27][3], c3[28][3]);
    csa a3_27_2 (s2[27][1], s2[27][0], c1[27][0], s3[27][2], c3[28][2]);
    csa a3_27_1 (c2[27][4], c2[27][3], c2[27][2], s3[27][1], c3[28][1]);
    csa a3_27_0 (c2[27][1], c2[27][0],      zero, s3[27][0], c3[28][0]);
    csa a3_26_3 (s2[26][4], s2[26][3], s2[26][2], s3[26][3], c3[27][3]);
    csa a3_26_2 (s2[26][1], s2[26][0], c1[26][0], s3[26][2], c3[27][2]);
    csa a3_26_1 (c2[26][4], c2[26][3], c2[26][2], s3[26][1], c3[27][1]);
    csa a3_26_0 (c2[26][1], c2[26][0],      zero, s3[26][0], c3[27][0]);
    csa a3_25_3 (s2[25][4], s2[25][3], s2[25][2], s3[25][3], c3[26][3]);
    csa a3_25_2 (s2[25][1], s2[25][0], c1[25][0], s3[25][2], c3[26][2]);
    csa a3_25_1 (c2[25][4], c2[25][3], c2[25][2], s3[25][1], c3[26][1]);
    csa a3_25_0 (c2[25][1], c2[25][0],      zero, s3[25][0], c3[26][0]);
    csa a3_24_3 (s2[24][4], s2[24][3], s2[24][2], s3[24][3], c3[25][3]);
    csa a3_24_2 (s2[24][1], s2[24][0], c1[24][0], s3[24][2], c3[25][2]);
    csa a3_24_1 (c2[24][4], c2[24][3], c2[24][2], s3[24][1], c3[25][1]);
    csa a3_24_0 (c2[24][1], c2[24][0],      zero, s3[24][0], c3[25][0]);
    csa a3_23_3 (s2[23][4], s2[23][3], s2[23][2], s3[23][3], c3[24][3]);
    csa a3_23_2 (s2[23][1], s2[23][0], c1[23][0], s3[23][2], c3[24][2]);
    csa a3_23_1 (c2[23][4], c2[23][3], c2[23][2], s3[23][1], c3[24][1]);
    csa a3_23_0 (c2[23][1], c2[23][0],      zero, s3[23][0], c3[24][0]);
    csa a3_22_2 (s2[22][4], s2[22][3], s2[22][2], s3[22][2], c3[23][2]);
    csa a3_22_1 (s2[22][1], s2[22][0], c2[22][4], s3[22][1], c3[23][1]);
    csa a3_22_0 (c2[22][3], c2[22][2], c2[22][1], s3[22][0], c3[23][0]);
    //     22:   c2[22][0]
    csa a3_21_2 (s2[21][4], s2[21][3], s2[21][2], s3[21][2], c3[22][2]);
    csa a3_21_1 (s2[21][1], s2[21][0], c2[21][4], s3[21][1], c3[22][1]);
    csa a3_21_0 (c2[21][3], c2[21][2], c2[21][1], s3[21][0], c3[22][0]);
    //     21:   c2[21][0]
    csa a3_20_2 (s2[20][4], s2[20][3], s2[20][2], s3[20][2], c3[21][2]);
    csa a3_20_1 (s2[20][1], s2[20][0], c2[20][3], s3[20][1], c3[21][1]);
    csa a3_20_0 (c2[20][2], c2[20][1], c2[20][0], s3[20][0], c3[21][0]);
    csa a3_19_2 (s2[19][3], s2[19][2], s2[19][1], s3[19][2], c3[20][2]);
    csa a3_19_1 (s2[19][0], c1[19][0], c2[19][3], s3[19][1], c3[20][1]);
    csa a3_19_0 (c2[19][2], c2[19][1], c2[19][0], s3[19][0], c3[20][0]);
    csa a3_18_2 (s2[18][3], s2[18][2], s2[18][1], s3[18][2], c3[19][2]);
    csa a3_18_1 (s2[18][0], c1[18][0], c2[18][3], s3[18][1], c3[19][1]);
    csa a3_18_0 (c2[18][2], c2[18][1], c2[18][0], s3[18][0], c3[19][0]);
    csa a3_17_2 (s2[17][3], s2[17][2], s2[17][1], s3[17][2], c3[18][2]);
    csa a3_17_1 (s2[17][0], c2[17][3], c2[17][2], s3[17][1], c3[18][1]);
    csa a3_17_0 (c2[17][1], c2[17][0],      zero, s3[17][0], c3[18][0]);
    csa a3_16_2 (s2[16][3], s2[16][2], s2[16][1], s3[16][2], c3[17][2]);
    csa a3_16_1 (s2[16][0], c2[16][3], c2[16][2], s3[16][1], c3[17][1]);
    csa a3_16_0 (c2[16][1], c2[16][0],      zero, s3[16][0], c3[17][0]);
    csa a3_15_1 (s2[15][3], s2[15][2], s2[15][1], s3[15][1], c3[16][1]);
    csa a3_15_0 (s2[15][0], c2[15][2], c2[15][1], s3[15][0], c3[16][0]);
    //     15:   c2[15][0]
    csa a3_14_1 (s2[14][2], s2[14][1], s2[14][0], s3[14][1], c3[15][1]);
    csa a3_14_0 (c1[14][0], c2[14][2], c2[14][1], s3[14][0], c3[15][0]);
    //     14:   c2[14][0]
    csa a3_13_1 (s2[13][2], s2[13][1], s2[13][0], s3[13][1], c3[14][1]);
    csa a3_13_0 (c2[13][2], c2[13][1], c2[13][0], s3[13][0], c3[14][0]);
    csa a3_12_1 (s2[12][2], s2[12][1], s2[12][0], s3[12][1], c3[13][1]);
    csa a3_12_0 (c2[12][2], c2[12][1], c2[12][0], s3[12][0], c3[13][0]);
    csa a3_11_1 (s2[11][2], s2[11][1], s2[11][0], s3[11][1], c3[12][1]);
    csa a3_11_0 (c2[11][1], c2[11][0],      zero, s3[11][0], c3[12][0]);
    csa a3_10_1 (s2[10][1], s2[10][0], c1[10][0], s3[10][1], c3[11][1]);
    csa a3_10_0 (c2[10][1], c2[10][0],      zero, s3[10][0], c3[11][0]);
    csa a3_09_1 (s2[09][1], s2[09][0], c1[09][0], s3[09][1], c3[10][1]);
    csa a3_09_0 (c2[09][1], c2[09][0],      zero, s3[09][0], c3[10][0]);
    csa a3_08_0 (s2[08][1], s2[08][0], c2[08][1], s3[08][0], c3[09][0]);
    //     08:   c2[08][0]
    csa a3_07_0 (s2[07][1], s2[07][0], c2[07][1], s3[07][0], c3[08][0]);
    //     07:   c2[07][0]
    csa a3_06_0 (s2[06][1], s2[06][0], c2[06][0], s3[06][0], c3[07][0]);
    csa a3_05_0 (s2[05][0], c1[05][0], c2[05][0], s3[05][0], c3[06][0]);
    csa a3_04_0 (s2[04][0], c2[04][0],      zero, s3[04][0], c3[05][0]);
    csa a3_03_0 (s2[03][0], c2[03][0],      zero, s3[03][0], c3[04][0]);
    //     02:   s2[02][0]
    //     01:   s1[01][0]
    //     00:   p[00][00]
    // level 4 ------------------------------------------------------------
    wire  [2:0] s4 [48:4];
    wire  [2:0] c4 [49:5];
    //     49:   c3[49][0]
    csa a4_48_0 (s3[48][0], c3[48][0],      zero, s4[48][0], c4[49][0]);
    csa a4_47_0 (s3[47][0], c3[47][0],      zero, s4[47][0], c4[48][0]);
    csa a4_46_0 (s3[46][0], c3[46][0],      zero, s4[46][0], c4[47][0]);
    csa a4_45_0 (s3[45][0], c3[45][0],      zero, s4[45][0], c4[46][0]);
    csa a4_44_0 (s3[44][0], c3[44][0],      zero, s4[44][0], c4[45][0]);
    csa a4_43_0 (s3[43][0], c2[43][0], c3[43][0], s4[43][0], c4[44][0]);
    csa a4_42_0 (s3[42][0], c2[42][0], c3[42][0], s4[42][0], c4[43][0]);
    csa a4_41_0 (s3[41][0], c2[41][0], c3[41][1], s4[41][0], c4[42][0]);
    //     41:   c3[41][0]
    csa a4_40_0 (s3[40][1], s3[40][0], c3[40][1], s4[40][0], c4[41][0]);
    //     40:   c3[40][0]
    csa a4_39_0 (s3[39][1], s3[39][0], c3[39][1], s4[39][0], c4[40][0]);
    //     39:   c3[39][0]
    csa a4_38_0 (s3[38][1], s3[38][0], c3[38][1], s4[38][0], c4[39][0]);
    //     38:   c3[38][0]
    csa a4_37_0 (s3[37][1], s3[37][0], c3[37][1], s4[37][0], c4[38][0]);
    //     37:   c3[37][0]
    csa a4_36_1 (s3[36][1], s3[36][0], c2[36][0], s4[36][1], c4[37][1]);
    csa a4_36_0 (c3[36][1], c3[36][0],      zero, s4[36][0], c4[37][0]);
    csa a4_35_1 (s3[35][1], s3[35][0], c2[35][0], s4[35][1], c4[36][1]);
    csa a4_35_0 (c3[35][2], c3[35][1], c3[35][0], s4[35][0], c4[36][0]);
    csa a4_34_1 (s3[34][2], s3[34][1], s3[34][0], s4[34][1], c4[35][1]);
    csa a4_34_0 (c3[34][2], c3[34][1], c3[34][0], s4[34][0], c4[35][0]);
    csa a4_33_1 (s3[33][2], s3[33][1], s3[33][0], s4[33][1], c4[34][1]);
    csa a4_33_0 (c3[33][2], c3[33][1], c3[33][0], s4[33][0], c4[34][0]);
    csa a4_32_1 (s3[32][2], s3[32][1], s3[32][0], s4[32][1], c4[33][1]);
    csa a4_32_0 (c3[32][2], c3[32][1], c3[32][0], s4[32][0], c4[33][0]);
    csa a4_31_1 (s3[31][2], s3[31][1], s3[31][0], s4[31][1], c4[32][1]);
    csa a4_31_0 (c3[31][2], c3[31][1], c3[31][0], s4[31][0], c4[32][0]);
    csa a4_30_1 (s3[30][2], s3[30][1], s3[30][0], s4[30][1], c4[31][1]);
    csa a4_30_0 (c2[30][0], c3[30][2], c3[30][1], s4[30][0], c4[31][0]);
    //     30:   c3[30][0]
    csa a4_29_1 (s3[29][2], s3[29][1], s3[29][0], s4[29][1], c4[30][1]);
    csa a4_29_0 (c2[29][0], c3[29][2], c3[29][1], s4[29][0], c4[30][0]);
    //     29:   c3[29][0]
    csa a4_28_2 (s3[28][2], s3[28][1], s3[28][0], s4[28][2], c4[29][2]);
    csa a4_28_1 (c2[28][0], c3[28][3], c3[28][2], s4[28][1], c4[29][1]);
    csa a4_28_0 (c3[28][1], c3[28][0],      zero, s4[28][0], c4[29][0]);
    csa a4_27_2 (s3[27][3], s3[27][2], s3[27][1], s4[27][2], c4[28][2]);
    csa a4_27_1 (s3[27][0], c3[27][3], c3[27][2], s4[27][1], c4[28][1]);
    csa a4_27_0 (c3[27][1], c3[27][0],      zero, s4[27][0], c4[28][0]);
    csa a4_26_2 (s3[26][3], s3[26][2], s3[26][1], s4[26][2], c4[27][2]);
    csa a4_26_1 (s3[26][0], c3[26][3], c3[26][2], s4[26][1], c4[27][1]);
    csa a4_26_0 (c3[26][1], c3[26][0],      zero, s4[26][0], c4[27][0]);
    csa a4_25_2 (s3[25][3], s3[25][2], s3[25][1], s4[25][2], c4[26][2]);
    csa a4_25_1 (s3[25][0], c3[25][3], c3[25][2], s4[25][1], c4[26][1]);
    csa a4_25_0 (c3[25][1], c3[25][0],      zero, s4[25][0], c4[26][0]);
    csa a4_24_2 (s3[24][3], s3[24][2], s3[24][1], s4[24][2], c4[25][2]);
    csa a4_24_1 (s3[24][0], c3[24][3], c3[24][2], s4[24][1], c4[25][1]);
    csa a4_24_0 (c3[24][1], c3[24][0],      zero, s4[24][0], c4[25][0]);
    csa a4_23_1 (s3[23][3], s3[23][2], s3[23][1], s4[23][1], c4[24][1]);
    csa a4_23_0 (s3[23][0], c3[23][2], c3[23][1], s4[23][0], c4[24][0]);
    //     23:   c3[23][0]
    csa a4_22_1 (s3[22][2], s3[22][1], s3[22][0], s4[22][1], c4[23][1]);
    csa a4_22_0 (c2[22][0], c3[22][2], c3[22][1], s4[22][0], c4[23][0]);
    //     22:   c3[22][0]
    csa a4_21_1 (s3[21][2], s3[21][1], s3[21][0], s4[21][1], c4[22][1]);
    csa a4_21_0 (c2[21][0], c3[21][2], c3[21][1], s4[21][0], c4[22][0]);
    //     21:   c3[21][0]
    csa a4_20_1 (s3[20][2], s3[20][1], s3[20][0], s4[20][1], c4[21][1]);
    csa a4_20_0 (c3[20][2], c3[20][1], c3[20][0], s4[20][0], c4[21][0]);
    csa a4_19_1 (s3[19][2], s3[19][1], s3[19][0], s4[19][1], c4[20][1]);
    csa a4_19_0 (c3[19][2], c3[19][1], c3[19][0], s4[19][0], c4[20][0]);
    csa a4_18_1 (s3[18][2], s3[18][1], s3[18][0], s4[18][1], c4[19][1]);
    csa a4_18_0 (c3[18][2], c3[18][1], c3[18][0], s4[18][0], c4[19][0]);
    csa a4_17_1 (s3[17][2], s3[17][1], s3[17][0], s4[17][1], c4[18][1]);
    csa a4_17_0 (c3[17][2], c3[17][1], c3[17][0], s4[17][0], c4[18][0]);
    csa a4_16_1 (s3[16][2], s3[16][1], s3[16][0], s4[16][1], c4[17][1]);
    csa a4_16_0 (c3[16][1], c3[16][0],      zero, s4[16][0], c4[17][0]);
    csa a4_15_1 (s3[15][1], s3[15][0], c2[15][0], s4[15][1], c4[16][1]);
    csa a4_15_0 (c3[15][1], c3[15][0],      zero, s4[15][0], c4[16][0]);
    csa a4_14_1 (s3[14][1], s3[14][0], c2[14][0], s4[14][1], c4[15][1]);
    csa a4_14_0 (c3[14][1], c3[14][0],      zero, s4[14][0], c4[15][0]);
    csa a4_13_0 (s3[13][1], s3[13][0], c3[13][1], s4[13][0], c4[14][0]);
    //     13:   c3[13][0]
    csa a4_12_0 (s3[12][1], s3[12][0], c3[12][1], s4[12][0], c4[13][0]);
    //     12:   c3[12][0]
    csa a4_11_0 (s3[11][1], s3[11][0], c3[11][1], s4[11][0], c4[12][0]);
    //     11:   c3[11][0]
    csa a4_10_0 (s3[10][1], s3[10][0], c3[10][1], s4[10][0], c4[11][0]);
    //     10:   c3[10][0]
    csa a4_09_0 (s3[09][1], s3[09][0], c3[09][0], s4[09][0], c4[10][0]);
    csa a4_08_0 (s3[08][0], c2[08][0], c3[08][0], s4[08][0], c4[09][0]);
    csa a4_07_0 (s3[07][0], c2[07][0], c3[07][0], s4[07][0], c4[08][0]);
    csa a4_06_0 (s3[06][0], c3[06][0],      zero, s4[06][0], c4[07][0]);
    csa a4_05_0 (s3[05][0], c3[05][0],      zero, s4[05][0], c4[06][0]);
    csa a4_04_0 (s3[04][0], c3[04][0],      zero, s4[04][0], c4[05][0]);
    //     03:   s3[03][0]
    //     02:   s2[02][0]
    //     01:   s1[01][0]
    //     00:   p[00][00]
    // level 5 ------------------------------------------------------------
    wire  [1:0] s5 [49:5];
    wire  [1:0] c5 [50:6];
    csa a5_49_0 (c3[49][0], c4[49][0],      zero, s5[49][0], c5[50][0]);
    csa a5_48_0 (s4[48][0], c4[48][0],      zero, s5[48][0], c5[49][0]);
    csa a5_47_0 (s4[47][0], c4[47][0],      zero, s5[47][0], c5[48][0]);
    csa a5_46_0 (s4[46][0], c4[46][0],      zero, s5[46][0], c5[47][0]);
    csa a5_45_0 (s4[45][0], c4[45][0],      zero, s5[45][0], c5[46][0]);
    csa a5_44_0 (s4[44][0], c4[44][0],      zero, s5[44][0], c5[45][0]);
    csa a5_43_0 (s4[43][0], c4[43][0],      zero, s5[43][0], c5[44][0]);
    csa a5_42_0 (s4[42][0], c4[42][0],      zero, s5[42][0], c5[43][0]);
    csa a5_41_0 (s4[41][0], c3[41][0], c4[41][0], s5[41][0], c5[42][0]);
    csa a5_40_0 (s4[40][0], c3[40][0], c4[40][0], s5[40][0], c5[41][0]);
    csa a5_39_0 (s4[39][0], c3[39][0], c4[39][0], s5[39][0], c5[40][0]);
    csa a5_38_0 (s4[38][0], c3[38][0], c4[38][0], s5[38][0], c5[39][0]);
    csa a5_37_0 (s4[37][0], c3[37][0], c4[37][1], s5[37][0], c5[38][0]);
    //     37:   c4[37][0]
    csa a5_36_0 (s4[36][1], s4[36][0], c4[36][1], s5[36][0], c5[37][0]);
    //     36:   c4[36][0]
    csa a5_35_0 (s4[35][1], s4[35][0], c4[35][1], s5[35][0], c5[36][0]);
    //     35:   c4[35][0]
    csa a5_34_0 (s4[34][1], s4[34][0], c4[34][1], s5[34][0], c5[35][0]);
    //     34:   c4[34][0]
    csa a5_33_0 (s4[33][1], s4[33][0], c4[33][1], s5[33][0], c5[34][0]);
    //     33:   c4[33][0]
    csa a5_32_0 (s4[32][1], s4[32][0], c4[32][1], s5[32][0], c5[33][0]);
    //     32:   c4[32][0]
    csa a5_31_0 (s4[31][1], s4[31][0], c4[31][1], s5[31][0], c5[32][0]);
    //     31:   c4[31][0]
    csa a5_30_1 (s4[30][1], s4[30][0], c3[30][0], s5[30][1], c5[31][1]);
    csa a5_30_0 (c4[30][1], c4[30][0],      zero, s5[30][0], c5[31][0]);
    csa a5_29_1 (s4[29][1], s4[29][0], c3[29][0], s5[29][1], c5[30][1]);
    csa a5_29_0 (c4[29][2], c4[29][1], c4[29][0], s5[29][0], c5[30][0]);
    csa a5_28_1 (s4[28][2], s4[28][1], s4[28][0], s5[28][1], c5[29][1]);
    csa a5_28_0 (c4[28][2], c4[28][1], c4[28][0], s5[28][0], c5[29][0]);
    csa a5_27_1 (s4[27][2], s4[27][1], s4[27][0], s5[27][1], c5[28][1]);
    csa a5_27_0 (c4[27][2], c4[27][1], c4[27][0], s5[27][0], c5[28][0]);
    csa a5_26_1 (s4[26][2], s4[26][1], s4[26][0], s5[26][1], c5[27][1]);
    csa a5_26_0 (c4[26][2], c4[26][1], c4[26][0], s5[26][0], c5[27][0]);
    csa a5_25_1 (s4[25][2], s4[25][1], s4[25][0], s5[25][1], c5[26][1]);
    csa a5_25_0 (c4[25][2], c4[25][1], c4[25][0], s5[25][0], c5[26][0]);
    csa a5_24_1 (s4[24][2], s4[24][1], s4[24][0], s5[24][1], c5[25][1]);
    csa a5_24_0 (c4[24][1], c4[24][0],      zero, s5[24][0], c5[25][0]);
    csa a5_23_1 (s4[23][1], s4[23][0], c3[23][0], s5[23][1], c5[24][1]);
    csa a5_23_0 (c4[23][1], c4[23][0],      zero, s5[23][0], c5[24][0]);
    csa a5_22_1 (s4[22][1], s4[22][0], c3[22][0], s5[22][1], c5[23][1]);
    csa a5_22_0 (c4[22][1], c4[22][0],      zero, s5[22][0], c5[23][0]);
    csa a5_21_1 (s4[21][1], s4[21][0], c3[21][0], s5[21][1], c5[22][1]);
    csa a5_21_0 (c4[21][1], c4[21][0],      zero, s5[21][0], c5[22][0]);
    csa a5_20_0 (s4[20][1], s4[20][0], c4[20][1], s5[20][0], c5[21][0]);
    //     20:   c4[20][0]
    csa a5_19_0 (s4[19][1], s4[19][0], c4[19][1], s5[19][0], c5[20][0]);
    //     19:   c4[19][0]
    csa a5_18_0 (s4[18][1], s4[18][0], c4[18][1], s5[18][0], c5[19][0]);
    //     18:   c4[18][0]
    csa a5_17_0 (s4[17][1], s4[17][0], c4[17][1], s5[17][0], c5[18][0]);
    //     17:   c4[17][0]
    csa a5_16_0 (s4[16][1], s4[16][0], c4[16][1], s5[16][0], c5[17][0]);
    //     16:   c4[16][0]
    csa a5_15_0 (s4[15][1], s4[15][0], c4[15][1], s5[15][0], c5[16][0]);
    //     15:   c4[15][0]
    csa a5_14_0 (s4[14][1], s4[14][0], c4[14][0], s5[14][0], c5[15][0]);
    csa a5_13_0 (s4[13][0], c3[13][0], c4[13][0], s5[13][0], c5[14][0]);
    csa a5_12_0 (s4[12][0], c3[12][0], c4[12][0], s5[12][0], c5[13][0]);
    csa a5_11_0 (s4[11][0], c3[11][0], c4[11][0], s5[11][0], c5[12][0]);
    csa a5_10_0 (s4[10][0], c3[10][0], c4[10][0], s5[10][0], c5[11][0]);
    csa a5_09_0 (s4[09][0], c4[09][0],      zero, s5[09][0], c5[10][0]);
    csa a5_08_0 (s4[08][0], c4[08][0],      zero, s5[08][0], c5[09][0]);
    csa a5_07_0 (s4[07][0], c4[07][0],      zero, s5[07][0], c5[08][0]);
    csa a5_06_0 (s4[06][0], c4[06][0],      zero, s5[06][0], c5[07][0]);
    csa a5_05_0 (s4[05][0], c4[05][0],      zero, s5[05][0], c5[06][0]);
    //     04:   s4[04][0]
    //     03:   s3[03][0]
    //     02:   s2[02][0]
    //     01:   s1[01][0]
    //     00:   p[00][00]
    // level 6 ------------------------------------------------------------
    wire  [0:0] s6 [49:6];
    wire  [0:0] c6 [50:7];
    csa a6_49_0 (s5[49][0], c5[49][0],      zero, s6[49][0], c6[50][0]);
    csa a6_48_0 (s5[48][0], c5[48][0],      zero, s6[48][0], c6[49][0]);
    csa a6_47_0 (s5[47][0], c5[47][0],      zero, s6[47][0], c6[48][0]);
    csa a6_46_0 (s5[46][0], c5[46][0],      zero, s6[46][0], c6[47][0]);
    csa a6_45_0 (s5[45][0], c5[45][0],      zero, s6[45][0], c6[46][0]);
    csa a6_44_0 (s5[44][0], c5[44][0],      zero, s6[44][0], c6[45][0]);
    csa a6_43_0 (s5[43][0], c5[43][0],      zero, s6[43][0], c6[44][0]);
    csa a6_42_0 (s5[42][0], c5[42][0],      zero, s6[42][0], c6[43][0]);
    csa a6_41_0 (s5[41][0], c5[41][0],      zero, s6[41][0], c6[42][0]);
    csa a6_40_0 (s5[40][0], c5[40][0],      zero, s6[40][0], c6[41][0]);
    csa a6_39_0 (s5[39][0], c5[39][0],      zero, s6[39][0], c6[40][0]);
    csa a6_38_0 (s5[38][0], c5[38][0],      zero, s6[38][0], c6[39][0]);
    csa a6_37_0 (s5[37][0], c4[37][0], c5[37][0], s6[37][0], c6[38][0]);
    csa a6_36_0 (s5[36][0], c4[36][0], c5[36][0], s6[36][0], c6[37][0]);
    csa a6_35_0 (s5[35][0], c4[35][0], c5[35][0], s6[35][0], c6[36][0]);
    csa a6_34_0 (s5[34][0], c4[34][0], c5[34][0], s6[34][0], c6[35][0]);
    csa a6_33_0 (s5[33][0], c4[33][0], c5[33][0], s6[33][0], c6[34][0]);
    csa a6_32_0 (s5[32][0], c4[32][0], c5[32][0], s6[32][0], c6[33][0]);
    csa a6_31_0 (s5[31][0], c4[31][0], c5[31][1], s6[31][0], c6[32][0]);
    //     31:   c5[31][0]
    csa a6_30_0 (s5[30][1], s5[30][0], c5[30][1], s6[30][0], c6[31][0]);
    //     30:   c5[30][0]
    csa a6_29_0 (s5[29][1], s5[29][0], c5[29][1], s6[29][0], c6[30][0]);
    //     29:   c5[29][0]
    csa a6_28_0 (s5[28][1], s5[28][0], c5[28][1], s6[28][0], c6[29][0]);
    //     28:   c5[28][0]
    csa a6_27_0 (s5[27][1], s5[27][0], c5[27][1], s6[27][0], c6[28][0]);
    //     27:   c5[27][0]
    csa a6_26_0 (s5[26][1], s5[26][0], c5[26][1], s6[26][0], c6[27][0]);
    //     26:   c5[26][0]
    csa a6_25_0 (s5[25][1], s5[25][0], c5[25][1], s6[25][0], c6[26][0]);
    //     25:   c5[25][0]
    csa a6_24_0 (s5[24][1], s5[24][0], c5[24][1], s6[24][0], c6[25][0]);
    //     24:   c5[24][0]
    csa a6_23_0 (s5[23][1], s5[23][0], c5[23][1], s6[23][0], c6[24][0]);
    //     23:   c5[23][0]
    csa a6_22_0 (s5[22][1], s5[22][0], c5[22][1], s6[22][0], c6[23][0]);
    //     22:   c5[22][0]
    csa a6_21_0 (s5[21][1], s5[21][0], c5[21][0], s6[21][0], c6[22][0]);
    csa a6_20_0 (s5[20][0], c4[20][0], c5[20][0], s6[20][0], c6[21][0]);
    csa a6_19_0 (s5[19][0], c4[19][0], c5[19][0], s6[19][0], c6[20][0]);
    csa a6_18_0 (s5[18][0], c4[18][0], c5[18][0], s6[18][0], c6[19][0]);
    csa a6_17_0 (s5[17][0], c4[17][0], c5[17][0], s6[17][0], c6[18][0]);
    csa a6_16_0 (s5[16][0], c4[16][0], c5[16][0], s6[16][0], c6[17][0]);
    csa a6_15_0 (s5[15][0], c4[15][0], c5[15][0], s6[15][0], c6[16][0]);
    csa a6_14_0 (s5[14][0], c5[14][0],      zero, s6[14][0], c6[15][0]);
    csa a6_13_0 (s5[13][0], c5[13][0],      zero, s6[13][0], c6[14][0]);
    csa a6_12_0 (s5[12][0], c5[12][0],      zero, s6[12][0], c6[13][0]);
    csa a6_11_0 (s5[11][0], c5[11][0],      zero, s6[11][0], c6[12][0]);
    csa a6_10_0 (s5[10][0], c5[10][0],      zero, s6[10][0], c6[11][0]);
    csa a6_09_0 (s5[09][0], c5[09][0],      zero, s6[09][0], c6[10][0]);
    csa a6_08_0 (s5[08][0], c5[08][0],      zero, s6[08][0], c6[09][0]);
    csa a6_07_0 (s5[07][0], c5[07][0],      zero, s6[07][0], c6[08][0]);
    csa a6_06_0 (s5[06][0], c5[06][0],      zero, s6[06][0], c6[07][0]);
    //     05:   s5[05][0]
    //     04:   s4[04][0]
    //     03:   s3[03][0]
    //     02:   s2[02][0]
    //     01:   s1[01][0]
    //     00:   p[00][00]
    // level 7 ------------------------------------------------------------
    wire  [0:0] s7 [49:7];
    wire  [0:0] c7 [50:8];
    csa a7_49_0 (s6[49][0], c6[49][0],      zero, s7[49][0], c7[50][0]);
    csa a7_48_0 (s6[48][0], c6[48][0],      zero, s7[48][0], c7[49][0]);
    csa a7_47_0 (s6[47][0], c6[47][0],      zero, s7[47][0], c7[48][0]);
    csa a7_46_0 (s6[46][0], c6[46][0],      zero, s7[46][0], c7[47][0]);
    csa a7_45_0 (s6[45][0], c6[45][0],      zero, s7[45][0], c7[46][0]);
    csa a7_44_0 (s6[44][0], c6[44][0],      zero, s7[44][0], c7[45][0]);
    csa a7_43_0 (s6[43][0], c6[43][0],      zero, s7[43][0], c7[44][0]);
    csa a7_42_0 (s6[42][0], c6[42][0],      zero, s7[42][0], c7[43][0]);
    csa a7_41_0 (s6[41][0], c6[41][0],      zero, s7[41][0], c7[42][0]);
    csa a7_40_0 (s6[40][0], c6[40][0],      zero, s7[40][0], c7[41][0]);
    csa a7_39_0 (s6[39][0], c6[39][0],      zero, s7[39][0], c7[40][0]);
    csa a7_38_0 (s6[38][0], c6[38][0],      zero, s7[38][0], c7[39][0]);
    csa a7_37_0 (s6[37][0], c6[37][0],      zero, s7[37][0], c7[38][0]);
    csa a7_36_0 (s6[36][0], c6[36][0],      zero, s7[36][0], c7[37][0]);
    csa a7_35_0 (s6[35][0], c6[35][0],      zero, s7[35][0], c7[36][0]);
    csa a7_34_0 (s6[34][0], c6[34][0],      zero, s7[34][0], c7[35][0]);
    csa a7_33_0 (s6[33][0], c6[33][0],      zero, s7[33][0], c7[34][0]);
    csa a7_32_0 (s6[32][0], c6[32][0],      zero, s7[32][0], c7[33][0]);
    csa a7_31_0 (s6[31][0], c5[31][0], c6[31][0], s7[31][0], c7[32][0]);
    csa a7_30_0 (s6[30][0], c5[30][0], c6[30][0], s7[30][0], c7[31][0]);
    csa a7_29_0 (s6[29][0], c5[29][0], c6[29][0], s7[29][0], c7[30][0]);
    csa a7_28_0 (s6[28][0], c5[28][0], c6[28][0], s7[28][0], c7[29][0]);
    csa a7_27_0 (s6[27][0], c5[27][0], c6[27][0], s7[27][0], c7[28][0]);
    csa a7_26_0 (s6[26][0], c5[26][0], c6[26][0], s7[26][0], c7[27][0]);
    csa a7_25_0 (s6[25][0], c5[25][0], c6[25][0], s7[25][0], c7[26][0]);
    csa a7_24_0 (s6[24][0], c5[24][0], c6[24][0], s7[24][0], c7[25][0]);
    csa a7_23_0 (s6[23][0], c5[23][0], c6[23][0], s7[23][0], c7[24][0]);
    csa a7_22_0 (s6[22][0], c5[22][0], c6[22][0], s7[22][0], c7[23][0]);
    csa a7_21_0 (s6[21][0], c6[21][0],      zero, s7[21][0], c7[22][0]);
    csa a7_20_0 (s6[20][0], c6[20][0],      zero, s7[20][0], c7[21][0]);
    csa a7_19_0 (s6[19][0], c6[19][0],      zero, s7[19][0], c7[20][0]);
    csa a7_18_0 (s6[18][0], c6[18][0],      zero, s7[18][0], c7[19][0]);
    csa a7_17_0 (s6[17][0], c6[17][0],      zero, s7[17][0], c7[18][0]);
    csa a7_16_0 (s6[16][0], c6[16][0],      zero, s7[16][0], c7[17][0]);
    csa a7_15_0 (s6[15][0], c6[15][0],      zero, s7[15][0], c7[16][0]);
    csa a7_14_0 (s6[14][0], c6[14][0],      zero, s7[14][0], c7[15][0]);
    csa a7_13_0 (s6[13][0], c6[13][0],      zero, s7[13][0], c7[14][0]);
    csa a7_12_0 (s6[12][0], c6[12][0],      zero, s7[12][0], c7[13][0]);
    csa a7_11_0 (s6[11][0], c6[11][0],      zero, s7[11][0], c7[12][0]);
    csa a7_10_0 (s6[10][0], c6[10][0],      zero, s7[10][0], c7[11][0]);
    csa a7_09_0 (s6[09][0], c6[09][0],      zero, s7[09][0], c7[10][0]);
    csa a7_08_0 (s6[08][0], c6[08][0],      zero, s7[08][0], c7[09][0]);
    csa a7_07_0 (s6[07][0], c6[07][0],      zero, s7[07][0], c7[08][0]);
    //     06:   s6[06][0]
    //     05:   s5[05][0]
    //     04:   s4[04][0]
    //     03:   s3[03][0]
    //     02:   s2[02][0]
    //     01:   s1[01][0]
    //     00:   p[00][00]
    assign x[49] = s7[49][0];                  assign y[49] = c7[49][0];
    assign x[48] = s7[48][0];                  assign y[48] = c7[48][0];
    assign x[47] = s7[47][0];                  assign y[47] = c7[47][0];
    assign x[46] = s7[46][0];                  assign y[46] = c7[46][0];
    assign x[45] = s7[45][0];                  assign y[45] = c7[45][0];
    assign x[44] = s7[44][0];                  assign y[44] = c7[44][0];
    assign x[43] = s7[43][0];                  assign y[43] = c7[43][0];
    assign x[42] = s7[42][0];                  assign y[42] = c7[42][0];
    assign x[41] = s7[41][0];                  assign y[41] = c7[41][0];
    assign x[40] = s7[40][0];                  assign y[40] = c7[40][0];
    assign x[39] = s7[39][0];                  assign y[39] = c7[39][0];
    assign x[38] = s7[38][0];                  assign y[38] = c7[38][0];
    assign x[37] = s7[37][0];                  assign y[37] = c7[37][0];
    assign x[36] = s7[36][0];                  assign y[36] = c7[36][0];
    assign x[35] = s7[35][0];                  assign y[35] = c7[35][0];
    assign x[34] = s7[34][0];                  assign y[34] = c7[34][0];
    assign x[33] = s7[33][0];                  assign y[33] = c7[33][0];
    assign x[32] = s7[32][0];                  assign y[32] = c7[32][0];
    assign x[31] = s7[31][0];                  assign y[31] = c7[31][0];
    assign x[30] = s7[30][0];                  assign y[30] = c7[30][0];
    assign x[29] = s7[29][0];                  assign y[29] = c7[29][0];
    assign x[28] = s7[28][0];                  assign y[28] = c7[28][0];
    assign x[27] = s7[27][0];                  assign y[27] = c7[27][0];
    assign x[26] = s7[26][0];                  assign y[26] = c7[26][0];
    assign x[25] = s7[25][0];                  assign y[25] = c7[25][0];
    assign x[24] = s7[24][0];                  assign y[24] = c7[24][0];
    assign x[23] = s7[23][0];                  assign y[23] = c7[23][0];
    assign x[22] = s7[22][0];                  assign y[22] = c7[22][0];
    assign x[21] = s7[21][0];                  assign y[21] = c7[21][0];
    assign x[20] = s7[20][0];                  assign y[20] = c7[20][0];
    assign x[19] = s7[19][0];                  assign y[19] = c7[19][0];
    assign x[18] = s7[18][0];                  assign y[18] = c7[18][0];
    assign x[17] = s7[17][0];                  assign y[17] = c7[17][0];
    assign x[16] = s7[16][0];                  assign y[16] = c7[16][0];
    assign x[15] = s7[15][0];                  assign y[15] = c7[15][0];
    assign x[14] = s7[14][0];                  assign y[14] = c7[14][0];
    assign x[13] = s7[13][0];                  assign y[13] = c7[13][0];
    assign x[12] = s7[12][0];                  assign y[12] = c7[12][0];
    assign x[11] = s7[11][0];                  assign y[11] = c7[11][0];
    assign x[10] = s7[10][0];                  assign y[10] = c7[10][0];
    assign x[09] = s7[09][0];                  assign y[09] = c7[09][0];
    assign x[08] = s7[08][0];                  assign y[08] = c7[08][0];
    assign z[07] = s7[07][0];
    assign z[06] = s6[06][0];
    assign z[05] = s5[05][0];
    assign z[04] = s4[04][0];
    assign z[03] = s3[03][0];
    assign z[02] = s2[02][0];
    assign z[01] = s1[01][0];
    assign z[00] = p[00][00];
endmodule
