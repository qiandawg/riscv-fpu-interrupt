`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/04/2017 12:12:07 PM
// Design Name: 
// Module Name: sccomp_sys
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

`include "mfp_ahb_const.vh"

module sc_interrupt_sys(
input                  SI_CLK100MHZ,
input                  lock,     
input                  SI_Reset_N,
input                   SI_ClkIn,
output [31:0]           inst,
output [31:0]           pc,
output [31:0]           aluout,
output [31:0]           memout,
input                   memclk,
input                   intr,
output                  inta,
input  [`MFP_N_SW-1 :0] IO_Switch,
input  [`MFP_N_PB-1 :0] IO_PB,
output [`MFP_N_LED-1:0] IO_LED,
output [ 7          :0] IO_7SEGEN_N,
output [ 6          :0] IO_7SEG_N,
output                  IO_BUZZ,                  
output                  IO_RGB_SPI_MOSI,
output                  IO_RGB_SPI_SCK,
output                  IO_RGB_SPI_CS,
output                  IO_RGB_DC,
output                  IO_RGB_RST,
output                  IO_RGB_VCC_EN,
output                  IO_RGB_PEN,
output                  IO_CS,
output                  IO_SCK,
input                   IO_SDO,
input                   UART_RX,
inout [4:1]             JB,
input [26:0]            counter);

wire[31:0] dataBus; //Currently driven data bus based on HSEL
wire[31:0] data_cpu; //data driven by cpu
wire[31:0] data_mem; //data driven by data memory
wire[31:0] data_gpio; //data driven by GPIO module


wire wmem;                           // write data memory
wire clk;
wire clrn;


wire dbg_resetn_cpu;
wire dbg_halt_cpu;

assign clk = SI_ClkIn;
assign clrn = SI_Reset_N & dbg_resetn_cpu;

// Qian added logic to fix timing issue due to high fanout for dbg_halt_cpu

// 2-FF sync (if dbg_halt_cpu is async to clk)
(* ASYNC_REG="TRUE", SHREG_EXTRACT="NO" *) reg halt_s0 = 1'b0;
(* ASYNC_REG="TRUE", SHREG_EXTRACT="NO" *) reg halt_s1 = 1'b0;
always @(posedge clk) begin
  halt_s0 <= dbg_halt_cpu;
  halt_s1 <= halt_s0;
end

// Replication-friendly buffer register
(* max_fanout = 64 *) reg halt_buf;
always @(posedge clk) begin
  halt_buf <= halt_s1;
end

//Qian logic add end


sccpu_intr cpu (
           clk, //Clock input
           clrn, //Reset input
           halt_buf, //Halt signal input generated by JTAG core
           halt_buf ? 32'b0 : inst, //Current instruction input from instruction memory (if CPU is halted, this is forced to 0/NOP)
           memout, //The IO/Data-Memory bus input data
           pc, //Output containing the current program counter (functions as the address on the instruction bus)
           wmem, //Output true when CPU is writing into IO/DMEM data bus
           aluout, //Output from ALU, drives the IO/DMEM address bus
           data_cpu, //Output containing the data to write into IO/DMEM data bus when wmem is true
           intr,
           int_sync,
           intr_ack  // interrupt acknowledge
           );
// Check if memory mapped I/O
wire[2:0] HSEL;


assign memout = dataBus;

//Be sure to use forward slashes '/', even on Windows
parameter IMEM_FILE = "C:/risc-fpu-interrupts/sc-interrupt/src/Assembly/RISCVscintSwitchLED7Seg/imem.mem";
parameter DMEM_FILE = "C:/risc-fpu-interrupts/sc-interrupt/src/Assembly/RISCVscintSwitchLED7Seg/dmem.mem";
//parameter IMEM_FILE = "C:/risc-fpu-interrupts/sc-interrupt/src/Assembly/RISCVsc_intTest/imem.mem";
//parameter DMEM_FILE = "C:/risc-fpu-interrupts/sc-interrupt/src/Assembly/RISCVsc_intTest/dmem.mem";

wire[31:0] dbg_imem_addr;
wire[31:0] dbg_imem_din;
wire dbg_imem_ce;
wire dbg_imem_we;

wire[31:0] dbg_dmem_addr;
wire[31:0] dbg_dmem_din;
wire dbg_dmem_ce;
wire dbg_dmem_we;

wire[31:0] effectiveIMemAddr = dbg_imem_ce ? dbg_imem_addr : pc;

uram #(.A_WIDTH(8), .INIT_FILE(IMEM_FILE), .READ_DELAY(0)) imem
    (.clk(clk), .we(dbg_imem_we), .cs(1'b1), .addr(effectiveIMemAddr), .data_in(dbg_imem_din), .data_out(inst));

wire effectiveDMemWE = dbg_dmem_ce ? dbg_dmem_we : wmem;
wire effectiveDMemCE = dbg_dmem_ce | HSEL[1];
wire[31:0] effectiveDMemAddr = dbg_dmem_ce ? dbg_dmem_addr : aluout;
uram #(.A_WIDTH(8), .INIT_FILE(DMEM_FILE), .READ_DELAY(0)) dmem
        (.clk(clk), .we(effectiveDMemWE), .cs(effectiveDMemCE), .addr(effectiveDMemAddr), .data_in(memout), .data_out(data_mem));
        
sccomp_decoder decode(aluout,HSEL);

cpugpio gpio (.clk(clk),
    .clrn(clrn),
    .dataout(data_gpio),
    .datain(memout),
    .haddr(aluout[7:2]),
    .we(wmem),
    .HSEL(HSEL[2]),
    .IO_Switch(IO_Switch),
    .IO_PB(IO_PB),
    .IO_LED(IO_LED),
    .IO_7SEGEN_N(IO_7SEGEN_N),
    .IO_7SEG_N(IO_7SEG_N),
    .IO_BUZZ(IO_BUZZ),                
    .IO_RGB_SPI_MOSI(IO_RGB_SPI_MOSI),
    .IO_RGB_SPI_SCK(IO_RGB_SPI_SCK),
    .IO_RGB_SPI_CS(IO_RGB_SPI_CS),
    .IO_RGB_DC(IO_RGB_DC),
    .IO_RGB_RST(IO_RGB_RST),
    .IO_RGB_VCC_EN(IO_RGB_VCC_EN),
    .IO_RGB_PEN(IO_RGB_PEN),
    .IO_SDO(IO_SDO),
    .IO_CS(IO_CS),
    .IO_SCK(IO_SCK));

    debug_control debug_if(.serial_tx(JB[2]), .serial_rx(JB[3]), .cpu_clk(clk),
        .sys_rstn(SI_Reset_N), .cpu_imem_addr(dbg_imem_addr), 
        .cpu_debug_to_imem_data(dbg_imem_din), .cpu_imem_to_debug_data(inst),
        .cpu_imem_we(dbg_imem_we), .cpu_imem_ce(dbg_imem_ce),
        .cpu_dmem_addr(dbg_dmem_addr), .cpu_debug_to_dmem_data(dbg_dmem_din),
        .cpu_imem_to_debug_data_ready(dbg_imem_ce & ~dbg_imem_we),
        .cpu_dmem_to_debug_data_ready(dbg_dmem_ce & ~dbg_dmem_we),
        .cpu_dmem_to_debug_data(data_mem), .cpu_dmem_we(dbg_dmem_we),
        .cpu_dmem_ce(dbg_dmem_ce), .cpu_resetn_cpu(dbg_resetn_cpu),
        .cpu_halt_cpu(dbg_halt_cpu));

assign dataBus = dbg_dmem_we ? dbg_dmem_din :
                wmem ? data_cpu :
                HSEL[1] ? data_mem :
                HSEL[2] ? data_gpio :
                32'b0;

//ila_0 my_ila (
//    .clk(SI_CLK100MHZ),                  // Clock used for ILA
//    .probe0(inst),          // Probe for data bus
//    .probe1(pc),       // Probe for address bus
//    .probe2(SI_ClkIn),   // Probe for control signal 1
//    .probe3(SI_Reset_N),    // Probe for control signal 2
//    .probe4(lock),
//    .probe5(counter),
//    .probe6(IO_Switch),
//    .probe7(IO_LED),
//    .probe8(dbg_imem_cs),
//    .probe9(dbg_imem_we),
//    .probe10(dbg_imem_addr),
//    .probe11(dbg_imem_din),
//    .probe12(dbg_dmem_cs),
//    .probe13(dbg_dmem_we),
//    .probe14(dbg_dmem_addr),
//    .probe15(dbg_dmem_din),
//    .probe16(dbg_halt_cpu),
//    .probe17(IO_7SEGEN_N),
//    .probe18(IO_7SEG_N),
//    .probe19(intr),    
//    .probe20(inta)
//    );

endmodule
